module display(state, HEX0);
    input logic [5:0] state;
    output logic [6:0] HEX0, HEX1;
    always_comb begin
        case (state)
                        // Light: 6543210`
            6'b000000: HEX0 = ~7'b0111111; // 0
            6'b000001: HEX0 = ~7'b0000110; // 1
            6'b000010: HEX0 = ~7'b1011011; // 2
            6'b000011: HEX0 = ~7'b1001111; // 3
            6'b000100: HEX0 = ~7'b1100110; // 4
            6'b000101: HEX0 = ~7'b1101101; // 5
            6'b000110: HEX0 = ~7'b1111101; // 6
            6'b000111: HEX0 = ~7'b0000111; // 7
            6'b001000: HEX0 = ~7'b1111111; // 8
            6'b001001: HEX0 = ~7'b1101111; // 9
            6'b001010: HEX0 = ~7'b0111111; // A
            6'b001011: HEX0 = ~7'b0000110; // B
            6'b001100: HEX0 = ~7'b1011011; // C
            6'b001101: HEX0 = ~7'b1001111; // D
            6'b001110: HEX0 = ~7'b1100110; // E
            6'b001111: HEX0 = ~7'b1101101; // F
            6'b010000: HEX0 = ~7'b1111101; // G
            6'b010001: HEX0 = ~7'b0000111; // H
            6'b010010: HEX0 = ~7'b1111111; // I
            6'b010011: HEX0 = ~7'b1101111; // J
            6'b010100: HEX0 = ~7'b0111111; // K
            6'b010101: HEX0 = ~7'b0000110; // L
            6'b010110: HEX0 = ~7'b1011011; // M
            6'b010111: HEX0 = ~7'b1001111; // N
            6'b011000: HEX0 = ~7'b1100110; // O
            6'b011001: HEX0 = ~7'b1101101; // P
            6'b011010: HEX0 = ~7'b1111101; // Q
            6'b011011: HEX0 = ~7'b0000111; // R
            6'b011100: HEX0 = ~7'b1111111; // S
            6'b011101: HEX0 = ~7'b1101111; // T
            6'b011110: HEX0 = ~7'b0111111; // U
            6'b011111: HEX0 = ~7'b0000110; // V
            6'b100000: HEX0 = ~7'b1011011; // W
            6'b100001: HEX0 = ~7'b1001111; // X
            6'b100010: HEX0 = ~7'b1100110; // Y
            6'b100011: HEX0 = ~7'b1101101; // Z
            6'b: HEX0 = ~7'b1111101; // special states 
            default:   
                begin
                       HEX0 = ~7'b1111111;
                       HEX1 = ~7'b1111111;
                end
        endcase
    end
endmodule